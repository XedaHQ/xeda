../blinky/ecp5pll.vhdl